module dummy();
    logic a;
    assign a = 1'b1;
endmodule
